// Gate-level modeling of NAND gate
module nand_gate (input a, input b, output y);
    nand (y, a, b); 
endmodule
