// Gate-level modeling of an AND gate
module and_gate (input a, input b, output y);
    and (y, a, b);
endmodule
